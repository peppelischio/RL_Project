------ Libraries and entity ------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

--- just two copied lines to start lol ---
